
package my_pkg;
`include "item.sv";
`include "Sequence.sv";
`include "Sequencer.sv";
`include "driver.sv";
`include "environment.sv";
`include "agent.sv";
`include "scoreboard.sv";
`include "monitor.sv";
`include "base_test.sv";
`include "func_cov.sv";
`include "testcase_1.sv";
`include "testcase_2.sv";
`include "testcase_3.sv";
`include "testcase_4.sv";
`include "testcase_5.sv";
`include "testcase_6.sv";
`include "testcase_7.sv";
`include "testcase_8.sv";
`include "testcase_9.sv";
`include "testcase_10.sv";
`include "testcase_11.sv";
`include "testcase_12.sv";
`include "testcase_13.sv";
`include "testcase_14.sv";
`include "testcase_15.sv";
`include "testcase_16.sv";
`include "testcase_17.sv";
endpackage

