`ifndef my_PKG_SV
`define my_PKG_SV

package my_pkg;
`include "item.sv";
`include "Sequence.sv";
`include "Sequencer.sv";
`include "driver.sv";
`include "environment.sv";
`include "agent.sv";
`include "scoreboard.sv";
`include "monitor.sv";
`include "base_test.sv";
`include "uvm_macros.svh";
endpackage
`endif
