interface add_if(input bit clk,reset);
  //logic reset;
  logic [3:0] ALU_Sel;
  logic [7:0] A;
  logic [7:0] B;
  logic [7:0] ALU_Out;
  logic CarryOut;

endinterface
